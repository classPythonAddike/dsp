`timescale 1ns/10ps

module DELAY_TB();
